package task_pkg;

  parameter [11:0] TASK_1_PKT_SIZE_IN_BYTES = 81;
  parameter [11:0] TASK_2_PKT_SIZE_IN_BYTES = 81;
  parameter [11:0] TASK_3_PKT_SIZE_IN_BYTES = 27;
  parameter [11:0] TASK_4_PKT_SIZE_IN_BYTES = 120;
  parameter [11:0] TASK_5_PKT_SIZE_IN_BYTES = 256;
  parameter [11:0] TASK_6_PKT_SIZE_IN_BYTES = 50;
  parameter [11:0] TASK_7_PKT_SIZE_IN_BYTES = 50;
  parameter [11:0] TASK_8_PKT_SIZE_IN_BYTES = 160;
  parameter [11:0] TASK_9_PKT_SIZE_IN_BYTES = 40;
  parameter [11:0] TASK_10_PKT_SIZE_IN_BYTES = 64;

endpackage 

