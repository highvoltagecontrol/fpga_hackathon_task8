//----------------------------------------------------------------------------------------
// TASK 9: 1/SQRT(X) 
// 
//----------------------------------------------------------------------------------------
module reciprocal_sqrt(i_clk, i_rst, i_enb, i_data, o_valid, o_data);

//-----		INPUTS		------------------------------------------------------------------	
		input i_clk;
		input i_rst;
		input i_enb;
		input [7:0] i_data;
//-----		OUTPUTS		------------------------------------------------------------------		
		output o_valid;
		output [31:0] o_data;
//-----    WIRES         -----------------------------------------------------------------
//-----    REGS         ------------------------------------------------------------------

//========================================================================================
//    		MODULE CONTENT		
//========================================================================================

		assign o_data = i_data; // Just a dummy assignement. Replace with your code.
		assign o_valid = i_enb; // Just a dummy assignement. Replace with your code.
		
endmodule 