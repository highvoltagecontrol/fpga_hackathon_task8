//----------------------------------------------------------------------------------------
// TASK 10: DEMODULATOR QAM16
// 
//----------------------------------------------------------------------------------------
module demod16(i_clk, i_data, i_rst, i_enb, o_data, o_valid);

//-----		INPUTS		----------------------------------------------------------	
	input i_clk;
	input [7:0] i_data;
	input i_rst;
	input i_enb;
//-----		OUTPUTS		----------------------------------------------------------		
	output [7:0] o_data;
	output o_valid;
//-----    WIRES         -----------------------------------------------------------------
//-----    REGS         ------------------------------------------------------------------
	
//========================================================================================
//    		MODULE CONTENT		
//========================================================================================

	assign o_data = i_data; // Just a dummy assignement. Replace with your code.
	assign o_valid = i_enb; // Just a dummy assignement. Replace with your code.
	
endmodule 